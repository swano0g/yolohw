`timescale 1ns / 1ps

module conv_pe #(
    parameter DATA_W = 8,
    parameter ACC_W  = 32
)(

);

endmodule
