`timescale 1ns / 1ps

module addr_sequencer;

parameter W_SIZE       = `W_SIZE;
parameter W_CHANNEL    = `W_CHANNEL;
parameter W_FRAME_SIZE = `W_FRAME_SIZE;
parameter Tin          = `Tin;
parameter Tout         = `Tout;

parameter IFM_AW       = `FM_BUFFER_AW;

parameter OFM_AW       = `FM_BUFFER_AW; 
localparam CLK_PERIOD       = 10; // 100 MHz


reg                  clk, rstn;
initial begin
    clk = 0; forever #(CLK_PERIOD/2) clk = ~clk;
end

reg  [W_SIZE-1:0]           q_width;
reg  [W_SIZE-1:0]           q_height;
reg  [W_CHANNEL-1:0]        q_channel;
reg  [W_CHANNEL-1:0]        q_channel_out;
reg  [W_SIZE+W_CHANNEL-1:0] q_row_stride;



//-------------------------------------------
// DUT: addr_sequencer
//-------------------------------------------
addr_sequencer u_addr_sequencer(
.clk(clk), 
.rstn(rstn),

// Addr Sequencer <-> TOP
.q_width(q_width),
.q_height(q_height),
.q_channel(q_channel),   
.q_channel_out(q_channel_out),
.q_row_stride(q_row_stride),   // q_width * q_channel


.q_addr_seq_start(),
.addr_seq_done(),

.q_as_mode(),          // 0 -> upsample, 1 -> route

.q_route_offset(),

// RD/WR addr 
.as_rd_vld(),
.as_rd_addr(),

// one cycle delay
.as_wr_vld(),
.as_wr_addr()
);

endmodule